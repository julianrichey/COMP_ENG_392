`timescale 1 ns / 1 ns

module softmax #(
    parameter integer DWIDTH_IN = 12, //8
    parameter integer DWIDTH_OUT = 12, //8
    parameter integer BITS = 10, //6
    parameter integer IMG_SIZE = 100
) (
    input clock,
    input reset,

    output reg fifo_in_rd_en,
    input [DWIDTH_IN-1:0] fifo_in_dout,
    input fifo_in_empty,
    output reg fifo_out_wr_en, 
    output reg [DWIDTH_OUT-1:0] fifo_out_din, 
    input fifo_out_full
);

localparam integer QUANT_VAL = 1 << BITS;
//localparam integer IMG_SIZE = 4096;//388800;

localparam integer BRAM_ADDR_WIDTH = 13;

reg [DWIDTH_OUT-1:0] fifo_out_din_c;
reg fifo_out_wr_en_c, bram_wr_en, move_on, move_on_c, move_on2, move_on2_c;

reg[BRAM_ADDR_WIDTH-1:0] bram_addr, bram_addr_c;

reg[DWIDTH_IN-1:0] bram_din, exp_val, exp_val_c;
wire[DWIDTH_IN-1:0] bram_dout;


integer denominator, denominator_c;
reg[DWIDTH_IN+BITS-1 : 0] alpha, alpha_c, mval; //converted_data

reg [2:0] state, next_state;
localparam PROLOGUE = 3'b000;
localparam MIDDLOGUE = 3'b001;
localparam BRAM_WR_STAGE = 3'b010;
localparam EPILOGUE = 3'b011;
localparam TEMP_END_STATE = 3'b100;

//reg my_in;

//reg[15:0] exp_arr[0:4095] = init_exp(my_in);
localparam[11:0] exp_arr [0:4096]= '{12'h012, 12'h012, 12'h012, 12'h012, 12'h012, 12'h012, 12'h012, 12'h012, 12'h012, 12'h012, 12'h012, 12'h012, 12'h012, 12'h012, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 
12'h013, 12'h013, 12'h013, 12'h013, 12'h013, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h014, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 12'h015, 
12'h015, 12'h015, 12'h015, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h016, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h017, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 
12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h018, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h019, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 
12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01a, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01b, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01c, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 
12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01d, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01e, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h01f, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 
12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h020, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h021, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h022, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 
12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h024, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h025, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h026, 12'h027, 12'h027, 12'h027, 12'h027, 12'h027, 12'h027, 12'h027, 12'h027, 12'h027, 12'h027, 12'h027, 
12'h027, 12'h027, 12'h027, 12'h027, 12'h027, 12'h027, 12'h027, 12'h027, 12'h027, 12'h027, 12'h027, 12'h027, 12'h027, 12'h027, 12'h027, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h028, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h029, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02a, 12'h02b, 12'h02b, 12'h02b, 12'h02b, 12'h02b, 12'h02b, 12'h02b, 12'h02b, 12'h02b, 12'h02b, 12'h02b, 
12'h02b, 12'h02b, 12'h02b, 12'h02b, 12'h02b, 12'h02b, 12'h02b, 12'h02b, 12'h02b, 12'h02b, 12'h02b, 12'h02b, 12'h02b, 12'h02c, 12'h02c, 12'h02c, 12'h02c, 12'h02c, 12'h02c, 12'h02c, 12'h02c, 12'h02c, 12'h02c, 12'h02c, 12'h02c, 12'h02c, 12'h02c, 12'h02c, 12'h02c, 12'h02c, 12'h02c, 12'h02c, 12'h02c, 12'h02c, 12'h02c, 12'h02c, 12'h02d, 12'h02d, 12'h02d, 12'h02d, 12'h02d, 12'h02d, 12'h02d, 12'h02d, 12'h02d, 12'h02d, 12'h02d, 12'h02d, 12'h02d, 12'h02d, 12'h02d, 12'h02d, 12'h02d, 12'h02d, 12'h02d, 12'h02d, 12'h02d, 12'h02d, 12'h02e, 12'h02e, 12'h02e, 12'h02e, 12'h02e, 12'h02e, 12'h02e, 12'h02e, 12'h02e, 12'h02e, 12'h02e, 12'h02e, 12'h02e, 12'h02e, 12'h02e, 12'h02e, 12'h02e, 12'h02e, 12'h02e, 12'h02e, 12'h02e, 12'h02e, 12'h02f, 12'h02f, 12'h02f, 12'h02f, 12'h02f, 12'h02f, 12'h02f, 12'h02f, 12'h02f, 12'h02f, 12'h02f, 12'h02f, 12'h02f, 12'h02f, 12'h02f, 12'h02f, 12'h02f, 12'h02f, 12'h02f, 12'h02f, 
12'h02f, 12'h02f, 12'h030, 12'h030, 12'h030, 12'h030, 12'h030, 12'h030, 12'h030, 12'h030, 12'h030, 12'h030, 12'h030, 12'h030, 12'h030, 12'h030, 12'h030, 12'h030, 12'h030, 12'h030, 12'h030, 12'h030, 12'h030, 12'h031, 12'h031, 12'h031, 12'h031, 12'h031, 12'h031, 12'h031, 12'h031, 12'h031, 12'h031, 12'h031, 12'h031, 12'h031, 12'h031, 12'h031, 12'h031, 12'h031, 12'h031, 12'h031, 12'h031, 12'h031, 12'h032, 12'h032, 12'h032, 12'h032, 12'h032, 12'h032, 12'h032, 12'h032, 12'h032, 12'h032, 12'h032, 12'h032, 12'h032, 12'h032, 12'h032, 12'h032, 12'h032, 12'h032, 12'h032, 12'h032, 12'h033, 12'h033, 12'h033, 12'h033, 12'h033, 12'h033, 12'h033, 12'h033, 12'h033, 12'h033, 12'h033, 12'h033, 12'h033, 12'h033, 12'h033, 12'h033, 12'h033, 12'h033, 12'h033, 12'h033, 12'h034, 12'h034, 12'h034, 12'h034, 12'h034, 12'h034, 12'h034, 12'h034, 12'h034, 12'h034, 12'h034, 12'h034, 12'h034, 12'h034, 12'h034, 12'h034, 
12'h034, 12'h034, 12'h034, 12'h035, 12'h035, 12'h035, 12'h035, 12'h035, 12'h035, 12'h035, 12'h035, 12'h035, 12'h035, 12'h035, 12'h035, 12'h035, 12'h035, 12'h035, 12'h035, 12'h035, 12'h035, 12'h035, 12'h036, 12'h036, 12'h036, 12'h036, 12'h036, 12'h036, 12'h036, 12'h036, 12'h036, 12'h036, 12'h036, 12'h036, 12'h036, 12'h036, 12'h036, 12'h036, 12'h036, 12'h036, 12'h036, 12'h037, 12'h037, 12'h037, 12'h037, 12'h037, 12'h037, 12'h037, 12'h037, 12'h037, 12'h037, 12'h037, 12'h037, 12'h037, 12'h037, 12'h037, 12'h037, 12'h037, 12'h037, 12'h037, 12'h038, 12'h038, 12'h038, 12'h038, 12'h038, 12'h038, 12'h038, 12'h038, 12'h038, 12'h038, 12'h038, 12'h038, 12'h038, 12'h038, 12'h038, 12'h038, 12'h038, 12'h038, 12'h039, 12'h039, 12'h039, 12'h039, 12'h039, 12'h039, 12'h039, 12'h039, 12'h039, 12'h039, 12'h039, 12'h039, 12'h039, 12'h039, 12'h039, 12'h039, 12'h039, 12'h039, 12'h03a, 12'h03a, 12'h03a, 12'h03a, 
12'h03a, 12'h03a, 12'h03a, 12'h03a, 12'h03a, 12'h03a, 12'h03a, 12'h03a, 12'h03a, 12'h03a, 12'h03a, 12'h03a, 12'h03a, 12'h03b, 12'h03b, 12'h03b, 12'h03b, 12'h03b, 12'h03b, 12'h03b, 12'h03b, 12'h03b, 12'h03b, 12'h03b, 12'h03b, 12'h03b, 12'h03b, 12'h03b, 12'h03b, 12'h03b, 12'h03c, 12'h03c, 12'h03c, 12'h03c, 12'h03c, 12'h03c, 12'h03c, 12'h03c, 12'h03c, 12'h03c, 12'h03c, 12'h03c, 12'h03c, 12'h03c, 12'h03c, 12'h03c, 12'h03c, 12'h03d, 12'h03d, 12'h03d, 12'h03d, 12'h03d, 12'h03d, 12'h03d, 12'h03d, 12'h03d, 12'h03d, 12'h03d, 12'h03d, 12'h03d, 12'h03d, 12'h03d, 12'h03d, 12'h03d, 12'h03e, 12'h03e, 12'h03e, 12'h03e, 12'h03e, 12'h03e, 12'h03e, 12'h03e, 12'h03e, 12'h03e, 12'h03e, 12'h03e, 12'h03e, 12'h03e, 12'h03e, 12'h03e, 12'h03f, 12'h03f, 12'h03f, 12'h03f, 12'h03f, 12'h03f, 12'h03f, 12'h03f, 12'h03f, 12'h03f, 12'h03f, 12'h03f, 12'h03f, 12'h03f, 12'h03f, 12'h03f, 12'h040, 12'h040, 12'h040, 12'h040, 
12'h040, 12'h040, 12'h040, 12'h040, 12'h040, 12'h040, 12'h040, 12'h040, 12'h040, 12'h040, 12'h040, 12'h040, 12'h041, 12'h041, 12'h041, 12'h041, 12'h041, 12'h041, 12'h041, 12'h041, 12'h041, 12'h041, 12'h041, 12'h041, 12'h041, 12'h041, 12'h041, 12'h041, 12'h042, 12'h042, 12'h042, 12'h042, 12'h042, 12'h042, 12'h042, 12'h042, 12'h042, 12'h042, 12'h042, 12'h042, 12'h042, 12'h042, 12'h042, 12'h043, 12'h043, 12'h043, 12'h043, 12'h043, 12'h043, 12'h043, 12'h043, 12'h043, 12'h043, 12'h043, 12'h043, 12'h043, 12'h043, 12'h043, 12'h044, 12'h044, 12'h044, 12'h044, 12'h044, 12'h044, 12'h044, 12'h044, 12'h044, 12'h044, 12'h044, 12'h044, 12'h044, 12'h044, 12'h044, 12'h045, 12'h045, 12'h045, 12'h045, 12'h045, 12'h045, 12'h045, 12'h045, 12'h045, 12'h045, 12'h045, 12'h045, 12'h045, 12'h045, 12'h045, 12'h046, 12'h046, 12'h046, 12'h046, 12'h046, 12'h046, 12'h046, 12'h046, 12'h046, 12'h046, 12'h046, 12'h046, 
12'h046, 12'h046, 12'h046, 12'h047, 12'h047, 12'h047, 12'h047, 12'h047, 12'h047, 12'h047, 12'h047, 12'h047, 12'h047, 12'h047, 12'h047, 12'h047, 12'h047, 12'h048, 12'h048, 12'h048, 12'h048, 12'h048, 12'h048, 12'h048, 12'h048, 12'h048, 12'h048, 12'h048, 12'h048, 12'h048, 12'h048, 12'h049, 12'h049, 12'h049, 12'h049, 12'h049, 12'h049, 12'h049, 12'h049, 12'h049, 12'h049, 12'h049, 12'h049, 12'h049, 12'h049, 12'h04a, 12'h04a, 12'h04a, 12'h04a, 12'h04a, 12'h04a, 12'h04a, 12'h04a, 12'h04a, 12'h04a, 12'h04a, 12'h04a, 12'h04a, 12'h04a, 12'h04b, 12'h04b, 12'h04b, 12'h04b, 12'h04b, 12'h04b, 12'h04b, 12'h04b, 12'h04b, 12'h04b, 12'h04b, 12'h04b, 12'h04b, 12'h04c, 12'h04c, 12'h04c, 12'h04c, 12'h04c, 12'h04c, 12'h04c, 12'h04c, 12'h04c, 12'h04c, 12'h04c, 12'h04c, 12'h04c, 12'h04c, 12'h04d, 12'h04d, 12'h04d, 12'h04d, 12'h04d, 12'h04d, 12'h04d, 12'h04d, 12'h04d, 12'h04d, 12'h04d, 12'h04d, 12'h04d, 12'h04e, 
12'h04e, 12'h04e, 12'h04e, 12'h04e, 12'h04e, 12'h04e, 12'h04e, 12'h04e, 12'h04e, 12'h04e, 12'h04e, 12'h04e, 12'h04f, 12'h04f, 12'h04f, 12'h04f, 12'h04f, 12'h04f, 12'h04f, 12'h04f, 12'h04f, 12'h04f, 12'h04f, 12'h04f, 12'h04f, 12'h050, 12'h050, 12'h050, 12'h050, 12'h050, 12'h050, 12'h050, 12'h050, 12'h050, 12'h050, 12'h050, 12'h050, 12'h050, 12'h051, 12'h051, 12'h051, 12'h051, 12'h051, 12'h051, 12'h051, 12'h051, 12'h051, 12'h051, 12'h051, 12'h051, 12'h052, 12'h052, 12'h052, 12'h052, 12'h052, 12'h052, 12'h052, 12'h052, 12'h052, 12'h052, 12'h052, 12'h052, 12'h052, 12'h053, 12'h053, 12'h053, 12'h053, 12'h053, 12'h053, 12'h053, 12'h053, 12'h053, 12'h053, 12'h053, 12'h053, 12'h054, 12'h054, 12'h054, 12'h054, 12'h054, 12'h054, 12'h054, 12'h054, 12'h054, 12'h054, 12'h054, 12'h054, 12'h055, 12'h055, 12'h055, 12'h055, 12'h055, 12'h055, 12'h055, 12'h055, 12'h055, 12'h055, 12'h055, 12'h055, 12'h056, 
12'h056, 12'h056, 12'h056, 12'h056, 12'h056, 12'h056, 12'h056, 12'h056, 12'h056, 12'h056, 12'h056, 12'h057, 12'h057, 12'h057, 12'h057, 12'h057, 12'h057, 12'h057, 12'h057, 12'h057, 12'h057, 12'h057, 12'h058, 12'h058, 12'h058, 12'h058, 12'h058, 12'h058, 12'h058, 12'h058, 12'h058, 12'h058, 12'h058, 12'h058, 12'h059, 12'h059, 12'h059, 12'h059, 12'h059, 12'h059, 12'h059, 12'h059, 12'h059, 12'h059, 12'h059, 12'h05a, 12'h05a, 12'h05a, 12'h05a, 12'h05a, 12'h05a, 12'h05a, 12'h05a, 12'h05a, 12'h05a, 12'h05a, 12'h05a, 12'h05b, 12'h05b, 12'h05b, 12'h05b, 12'h05b, 12'h05b, 12'h05b, 12'h05b, 12'h05b, 12'h05b, 12'h05b, 12'h05c, 12'h05c, 12'h05c, 12'h05c, 12'h05c, 12'h05c, 12'h05c, 12'h05c, 12'h05c, 12'h05c, 12'h05c, 12'h05d, 12'h05d, 12'h05d, 12'h05d, 12'h05d, 12'h05d, 12'h05d, 12'h05d, 12'h05d, 12'h05d, 12'h05d, 12'h05e, 12'h05e, 12'h05e, 12'h05e, 12'h05e, 12'h05e, 12'h05e, 12'h05e, 12'h05e, 12'h05e, 
12'h05e, 12'h05f, 12'h05f, 12'h05f, 12'h05f, 12'h05f, 12'h05f, 12'h05f, 12'h05f, 12'h05f, 12'h05f, 12'h05f, 12'h060, 12'h060, 12'h060, 12'h060, 12'h060, 12'h060, 12'h060, 12'h060, 12'h060, 12'h060, 12'h061, 12'h061, 12'h061, 12'h061, 12'h061, 12'h061, 12'h061, 12'h061, 12'h061, 12'h061, 12'h061, 12'h062, 12'h062, 12'h062, 12'h062, 12'h062, 12'h062, 12'h062, 12'h062, 12'h062, 12'h062, 12'h063, 12'h063, 12'h063, 12'h063, 12'h063, 12'h063, 12'h063, 12'h063, 12'h063, 12'h063, 12'h064, 12'h064, 12'h064, 12'h064, 12'h064, 12'h064, 12'h064, 12'h064, 12'h064, 12'h064, 12'h064, 12'h065, 12'h065, 12'h065, 12'h065, 12'h065, 12'h065, 12'h065, 12'h065, 12'h065, 12'h065, 12'h066, 12'h066, 12'h066, 12'h066, 12'h066, 12'h066, 12'h066, 12'h066, 12'h066, 12'h066, 12'h067, 12'h067, 12'h067, 12'h067, 12'h067, 12'h067, 12'h067, 12'h067, 12'h067, 12'h067, 12'h068, 12'h068, 12'h068, 12'h068, 12'h068, 12'h068, 
12'h068, 12'h068, 12'h068, 12'h069, 12'h069, 12'h069, 12'h069, 12'h069, 12'h069, 12'h069, 12'h069, 12'h069, 12'h069, 12'h06a, 12'h06a, 12'h06a, 12'h06a, 12'h06a, 12'h06a, 12'h06a, 12'h06a, 12'h06a, 12'h06a, 12'h06b, 12'h06b, 12'h06b, 12'h06b, 12'h06b, 12'h06b, 12'h06b, 12'h06b, 12'h06b, 12'h06c, 12'h06c, 12'h06c, 12'h06c, 12'h06c, 12'h06c, 12'h06c, 12'h06c, 12'h06c, 12'h06c, 12'h06d, 12'h06d, 12'h06d, 12'h06d, 12'h06d, 12'h06d, 12'h06d, 12'h06d, 12'h06d, 12'h06e, 12'h06e, 12'h06e, 12'h06e, 12'h06e, 12'h06e, 12'h06e, 12'h06e, 12'h06e, 12'h06f, 12'h06f, 12'h06f, 12'h06f, 12'h06f, 12'h06f, 12'h06f, 12'h06f, 12'h06f, 12'h070, 12'h070, 12'h070, 12'h070, 12'h070, 12'h070, 12'h070, 12'h070, 12'h070, 12'h070, 12'h071, 12'h071, 12'h071, 12'h071, 12'h071, 12'h071, 12'h071, 12'h071, 12'h071, 12'h072, 12'h072, 12'h072, 12'h072, 12'h072, 12'h072, 12'h072, 12'h072, 12'h073, 12'h073, 12'h073, 12'h073, 
12'h073, 12'h073, 12'h073, 12'h073, 12'h073, 12'h074, 12'h074, 12'h074, 12'h074, 12'h074, 12'h074, 12'h074, 12'h074, 12'h074, 12'h075, 12'h075, 12'h075, 12'h075, 12'h075, 12'h075, 12'h075, 12'h075, 12'h075, 12'h076, 12'h076, 12'h076, 12'h076, 12'h076, 12'h076, 12'h076, 12'h076, 12'h077, 12'h077, 12'h077, 12'h077, 12'h077, 12'h077, 12'h077, 12'h077, 12'h077, 12'h078, 12'h078, 12'h078, 12'h078, 12'h078, 12'h078, 12'h078, 12'h078, 12'h078, 12'h079, 12'h079, 12'h079, 12'h079, 12'h079, 12'h079, 12'h079, 12'h079, 12'h07a, 12'h07a, 12'h07a, 12'h07a, 12'h07a, 12'h07a, 12'h07a, 12'h07a, 12'h07b, 12'h07b, 12'h07b, 12'h07b, 12'h07b, 12'h07b, 12'h07b, 12'h07b, 12'h07b, 12'h07c, 12'h07c, 12'h07c, 12'h07c, 12'h07c, 12'h07c, 12'h07c, 12'h07c, 12'h07d, 12'h07d, 12'h07d, 12'h07d, 12'h07d, 12'h07d, 12'h07d, 12'h07d, 12'h07e, 12'h07e, 12'h07e, 12'h07e, 12'h07e, 12'h07e, 12'h07e, 12'h07e, 12'h07f, 12'h07f, 
12'h07f, 12'h07f, 12'h07f, 12'h07f, 12'h07f, 12'h07f, 12'h080, 12'h080, 12'h080, 12'h080, 12'h080, 12'h080, 12'h080, 12'h080, 12'h081, 12'h081, 12'h081, 12'h081, 12'h081, 12'h081, 12'h081, 12'h081, 12'h082, 12'h082, 12'h082, 12'h082, 12'h082, 12'h082, 12'h082, 12'h082, 12'h083, 12'h083, 12'h083, 12'h083, 12'h083, 12'h083, 12'h083, 12'h083, 12'h084, 12'h084, 12'h084, 12'h084, 12'h084, 12'h084, 12'h084, 12'h085, 12'h085, 12'h085, 12'h085, 12'h085, 12'h085, 12'h085, 12'h085, 12'h086, 12'h086, 12'h086, 12'h086, 12'h086, 12'h086, 12'h086, 12'h086, 12'h087, 12'h087, 12'h087, 12'h087, 12'h087, 12'h087, 12'h087, 12'h088, 12'h088, 12'h088, 12'h088, 12'h088, 12'h088, 12'h088, 12'h088, 12'h089, 12'h089, 12'h089, 12'h089, 12'h089, 12'h089, 12'h089, 12'h08a, 12'h08a, 12'h08a, 12'h08a, 12'h08a, 12'h08a, 12'h08a, 12'h08a, 12'h08b, 12'h08b, 12'h08b, 12'h08b, 12'h08b, 12'h08b, 12'h08b, 12'h08c, 12'h08c, 
12'h08c, 12'h08c, 12'h08c, 12'h08c, 12'h08c, 12'h08d, 12'h08d, 12'h08d, 12'h08d, 12'h08d, 12'h08d, 12'h08d, 12'h08e, 12'h08e, 12'h08e, 12'h08e, 12'h08e, 12'h08e, 12'h08e, 12'h08e, 12'h08f, 12'h08f, 12'h08f, 12'h08f, 12'h08f, 12'h08f, 12'h08f, 12'h090, 12'h090, 12'h090, 12'h090, 12'h090, 12'h090, 12'h090, 12'h091, 12'h091, 12'h091, 12'h091, 12'h091, 12'h091, 12'h091, 12'h092, 12'h092, 12'h092, 12'h092, 12'h092, 12'h092, 12'h092, 12'h093, 12'h093, 12'h093, 12'h093, 12'h093, 12'h093, 12'h093, 12'h094, 12'h094, 12'h094, 12'h094, 12'h094, 12'h094, 12'h094, 12'h095, 12'h095, 12'h095, 12'h095, 12'h095, 12'h095, 12'h095, 12'h096, 12'h096, 12'h096, 12'h096, 12'h096, 12'h096, 12'h097, 12'h097, 12'h097, 12'h097, 12'h097, 12'h097, 12'h097, 12'h098, 12'h098, 12'h098, 12'h098, 12'h098, 12'h098, 12'h098, 12'h099, 12'h099, 12'h099, 12'h099, 12'h099, 12'h099, 12'h099, 12'h09a, 12'h09a, 12'h09a, 12'h09a, 
12'h09a, 12'h09a, 12'h09b, 12'h09b, 12'h09b, 12'h09b, 12'h09b, 12'h09b, 12'h09b, 12'h09c, 12'h09c, 12'h09c, 12'h09c, 12'h09c, 12'h09c, 12'h09d, 12'h09d, 12'h09d, 12'h09d, 12'h09d, 12'h09d, 12'h09d, 12'h09e, 12'h09e, 12'h09e, 12'h09e, 12'h09e, 12'h09e, 12'h09f, 12'h09f, 12'h09f, 12'h09f, 12'h09f, 12'h09f, 12'h09f, 12'h0a0, 12'h0a0, 12'h0a0, 12'h0a0, 12'h0a0, 12'h0a0, 12'h0a1, 12'h0a1, 12'h0a1, 12'h0a1, 12'h0a1, 12'h0a1, 12'h0a2, 12'h0a2, 12'h0a2, 12'h0a2, 12'h0a2, 12'h0a2, 12'h0a2, 12'h0a3, 12'h0a3, 12'h0a3, 12'h0a3, 12'h0a3, 12'h0a3, 12'h0a4, 12'h0a4, 12'h0a4, 12'h0a4, 12'h0a4, 12'h0a4, 12'h0a5, 12'h0a5, 12'h0a5, 12'h0a5, 12'h0a5, 12'h0a5, 12'h0a6, 12'h0a6, 12'h0a6, 12'h0a6, 12'h0a6, 12'h0a6, 12'h0a7, 12'h0a7, 12'h0a7, 12'h0a7, 12'h0a7, 12'h0a7, 12'h0a7, 12'h0a8, 12'h0a8, 12'h0a8, 12'h0a8, 12'h0a8, 12'h0a8, 12'h0a9, 12'h0a9, 12'h0a9, 12'h0a9, 12'h0a9, 12'h0a9, 12'h0aa, 12'h0aa, 12'h0aa, 
12'h0aa, 12'h0aa, 12'h0aa, 12'h0ab, 12'h0ab, 12'h0ab, 12'h0ab, 12'h0ab, 12'h0ab, 12'h0ac, 12'h0ac, 12'h0ac, 12'h0ac, 12'h0ac, 12'h0ac, 12'h0ad, 12'h0ad, 12'h0ad, 12'h0ad, 12'h0ad, 12'h0ad, 12'h0ae, 12'h0ae, 12'h0ae, 12'h0ae, 12'h0ae, 12'h0af, 12'h0af, 12'h0af, 12'h0af, 12'h0af, 12'h0af, 12'h0b0, 12'h0b0, 12'h0b0, 12'h0b0, 12'h0b0, 12'h0b0, 12'h0b1, 12'h0b1, 12'h0b1, 12'h0b1, 12'h0b1, 12'h0b1, 12'h0b2, 12'h0b2, 12'h0b2, 12'h0b2, 12'h0b2, 12'h0b2, 12'h0b3, 12'h0b3, 12'h0b3, 12'h0b3, 12'h0b3, 12'h0b4, 12'h0b4, 12'h0b4, 12'h0b4, 12'h0b4, 12'h0b4, 12'h0b5, 12'h0b5, 12'h0b5, 12'h0b5, 12'h0b5, 12'h0b5, 12'h0b6, 12'h0b6, 12'h0b6, 12'h0b6, 12'h0b6, 12'h0b7, 12'h0b7, 12'h0b7, 12'h0b7, 12'h0b7, 12'h0b7, 12'h0b8, 12'h0b8, 12'h0b8, 12'h0b8, 12'h0b8, 12'h0b9, 12'h0b9, 12'h0b9, 12'h0b9, 12'h0b9, 12'h0b9, 12'h0ba, 12'h0ba, 12'h0ba, 12'h0ba, 12'h0ba, 12'h0bb, 12'h0bb, 12'h0bb, 12'h0bb, 12'h0bb, 12'h0bb, 
12'h0bc, 12'h0bc, 12'h0bc, 12'h0bc, 12'h0bc, 12'h0bd, 12'h0bd, 12'h0bd, 12'h0bd, 12'h0bd, 12'h0bd, 12'h0be, 12'h0be, 12'h0be, 12'h0be, 12'h0be, 12'h0bf, 12'h0bf, 12'h0bf, 12'h0bf, 12'h0bf, 12'h0c0, 12'h0c0, 12'h0c0, 12'h0c0, 12'h0c0, 12'h0c0, 12'h0c1, 12'h0c1, 12'h0c1, 12'h0c1, 12'h0c1, 12'h0c2, 12'h0c2, 12'h0c2, 12'h0c2, 12'h0c2, 12'h0c3, 12'h0c3, 12'h0c3, 12'h0c3, 12'h0c3, 12'h0c4, 12'h0c4, 12'h0c4, 12'h0c4, 12'h0c4, 12'h0c4, 12'h0c5, 12'h0c5, 12'h0c5, 12'h0c5, 12'h0c5, 12'h0c6, 12'h0c6, 12'h0c6, 12'h0c6, 12'h0c6, 12'h0c7, 12'h0c7, 12'h0c7, 12'h0c7, 12'h0c7, 12'h0c8, 12'h0c8, 12'h0c8, 12'h0c8, 12'h0c8, 12'h0c9, 12'h0c9, 12'h0c9, 12'h0c9, 12'h0c9, 12'h0ca, 12'h0ca, 12'h0ca, 12'h0ca, 12'h0ca, 12'h0cb, 12'h0cb, 12'h0cb, 12'h0cb, 12'h0cb, 12'h0cc, 12'h0cc, 12'h0cc, 12'h0cc, 12'h0cc, 12'h0cd, 12'h0cd, 12'h0cd, 12'h0cd, 12'h0cd, 12'h0ce, 12'h0ce, 12'h0ce, 12'h0ce, 12'h0ce, 12'h0cf, 12'h0cf, 
12'h0cf, 12'h0cf, 12'h0cf, 12'h0d0, 12'h0d0, 12'h0d0, 12'h0d0, 12'h0d0, 12'h0d1, 12'h0d1, 12'h0d1, 12'h0d1, 12'h0d1, 12'h0d2, 12'h0d2, 12'h0d2, 12'h0d2, 12'h0d2, 12'h0d3, 12'h0d3, 12'h0d3, 12'h0d3, 12'h0d3, 12'h0d4, 12'h0d4, 12'h0d4, 12'h0d4, 12'h0d4, 12'h0d5, 12'h0d5, 12'h0d5, 12'h0d5, 12'h0d6, 12'h0d6, 12'h0d6, 12'h0d6, 12'h0d6, 12'h0d7, 12'h0d7, 12'h0d7, 12'h0d7, 12'h0d7, 12'h0d8, 12'h0d8, 12'h0d8, 12'h0d8, 12'h0d8, 12'h0d9, 12'h0d9, 12'h0d9, 12'h0d9, 12'h0da, 12'h0da, 12'h0da, 12'h0da, 12'h0da, 12'h0db, 12'h0db, 12'h0db, 12'h0db, 12'h0db, 12'h0dc, 12'h0dc, 12'h0dc, 12'h0dc, 12'h0dd, 12'h0dd, 12'h0dd, 12'h0dd, 12'h0dd, 12'h0de, 12'h0de, 12'h0de, 12'h0de, 12'h0de, 12'h0df, 12'h0df, 12'h0df, 12'h0df, 12'h0e0, 12'h0e0, 12'h0e0, 12'h0e0, 12'h0e0, 12'h0e1, 12'h0e1, 12'h0e1, 12'h0e1, 12'h0e2, 12'h0e2, 12'h0e2, 12'h0e2, 12'h0e2, 12'h0e3, 12'h0e3, 12'h0e3, 12'h0e3, 12'h0e4, 12'h0e4, 12'h0e4, 
12'h0e4, 12'h0e4, 12'h0e5, 12'h0e5, 12'h0e5, 12'h0e5, 12'h0e6, 12'h0e6, 12'h0e6, 12'h0e6, 12'h0e6, 12'h0e7, 12'h0e7, 12'h0e7, 12'h0e7, 12'h0e8, 12'h0e8, 12'h0e8, 12'h0e8, 12'h0e8, 12'h0e9, 12'h0e9, 12'h0e9, 12'h0e9, 12'h0ea, 12'h0ea, 12'h0ea, 12'h0ea, 12'h0eb, 12'h0eb, 12'h0eb, 12'h0eb, 12'h0eb, 12'h0ec, 12'h0ec, 12'h0ec, 12'h0ec, 12'h0ed, 12'h0ed, 12'h0ed, 12'h0ed, 12'h0ee, 12'h0ee, 12'h0ee, 12'h0ee, 12'h0ee, 12'h0ef, 12'h0ef, 12'h0ef, 12'h0ef, 12'h0f0, 12'h0f0, 12'h0f0, 12'h0f0, 12'h0f1, 12'h0f1, 12'h0f1, 12'h0f1, 12'h0f2, 12'h0f2, 12'h0f2, 12'h0f2, 12'h0f2, 12'h0f3, 12'h0f3, 12'h0f3, 12'h0f3, 12'h0f4, 12'h0f4, 12'h0f4, 12'h0f4, 12'h0f5, 12'h0f5, 12'h0f5, 12'h0f5, 12'h0f6, 12'h0f6, 12'h0f6, 12'h0f6, 12'h0f7, 12'h0f7, 12'h0f7, 12'h0f7, 12'h0f8, 12'h0f8, 12'h0f8, 12'h0f8, 12'h0f8, 12'h0f9, 12'h0f9, 12'h0f9, 12'h0f9, 12'h0fa, 12'h0fa, 12'h0fa, 12'h0fa, 12'h0fb, 12'h0fb, 12'h0fb, 12'h0fb, 
12'h0fc, 12'h0fc, 12'h0fc, 12'h0fc, 12'h0fd, 12'h0fd, 12'h0fd, 12'h0fd, 12'h0fe, 12'h0fe, 12'h0fe, 12'h0fe, 12'h0ff, 12'h0ff, 12'h0ff, 12'h0ff, 12'h100, 12'h100, 12'h100, 12'h100, 12'h101, 12'h101, 12'h101, 12'h101, 12'h102, 12'h102, 12'h102, 12'h102, 12'h103, 12'h103, 12'h103, 12'h103, 12'h104, 12'h104, 12'h104, 12'h104, 12'h105, 12'h105, 12'h105, 12'h105, 12'h106, 12'h106, 12'h106, 12'h106, 12'h107, 12'h107, 12'h107, 12'h108, 12'h108, 12'h108, 12'h108, 12'h109, 12'h109, 12'h109, 12'h109, 12'h10a, 12'h10a, 12'h10a, 12'h10a, 12'h10b, 12'h10b, 12'h10b, 12'h10b, 12'h10c, 12'h10c, 12'h10c, 12'h10c, 12'h10d, 12'h10d, 12'h10d, 12'h10e, 12'h10e, 12'h10e, 12'h10e, 12'h10f, 12'h10f, 12'h10f, 12'h10f, 12'h110, 12'h110, 12'h110, 12'h110, 12'h111, 12'h111, 12'h111, 12'h111, 12'h112, 12'h112, 12'h112, 12'h113, 12'h113, 12'h113, 12'h113, 12'h114, 12'h114, 12'h114, 12'h114, 12'h115, 12'h115, 12'h115, 
12'h116, 12'h116, 12'h116, 12'h116, 12'h117, 12'h117, 12'h117, 12'h117, 12'h118, 12'h118, 12'h118, 12'h119, 12'h119, 12'h119, 12'h119, 12'h11a, 12'h11a, 12'h11a, 12'h11a, 12'h11b, 12'h11b, 12'h11b, 12'h11c, 12'h11c, 12'h11c, 12'h11c, 12'h11d, 12'h11d, 12'h11d, 12'h11e, 12'h11e, 12'h11e, 12'h11e, 12'h11f, 12'h11f, 12'h11f, 12'h11f, 12'h120, 12'h120, 12'h120, 12'h121, 12'h121, 12'h121, 12'h121, 12'h122, 12'h122, 12'h122, 12'h123, 12'h123, 12'h123, 12'h123, 12'h124, 12'h124, 12'h124, 12'h125, 12'h125, 12'h125, 12'h125, 12'h126, 12'h126, 12'h126, 12'h127, 12'h127, 12'h127, 12'h127, 12'h128, 12'h128, 12'h128, 12'h129, 12'h129, 12'h129, 12'h12a, 12'h12a, 12'h12a, 12'h12a, 12'h12b, 12'h12b, 12'h12b, 12'h12c, 12'h12c, 12'h12c, 12'h12c, 12'h12d, 12'h12d, 12'h12d, 12'h12e, 12'h12e, 12'h12e, 12'h12e, 12'h12f, 12'h12f, 12'h12f, 12'h130, 12'h130, 12'h130, 12'h131, 12'h131, 12'h131, 12'h131, 12'h132, 
12'h132, 12'h132, 12'h133, 12'h133, 12'h133, 12'h134, 12'h134, 12'h134, 12'h134, 12'h135, 12'h135, 12'h135, 12'h136, 12'h136, 12'h136, 12'h137, 12'h137, 12'h137, 12'h137, 12'h138, 12'h138, 12'h138, 12'h139, 12'h139, 12'h139, 12'h13a, 12'h13a, 12'h13a, 12'h13b, 12'h13b, 12'h13b, 12'h13b, 12'h13c, 12'h13c, 12'h13c, 12'h13d, 12'h13d, 12'h13d, 12'h13e, 12'h13e, 12'h13e, 12'h13f, 12'h13f, 12'h13f, 12'h140, 12'h140, 12'h140, 12'h140, 12'h141, 12'h141, 12'h141, 12'h142, 12'h142, 12'h142, 12'h143, 12'h143, 12'h143, 12'h144, 12'h144, 12'h144, 12'h145, 12'h145, 12'h145, 12'h146, 12'h146, 12'h146, 12'h146, 12'h147, 12'h147, 12'h147, 12'h148, 12'h148, 12'h148, 12'h149, 12'h149, 12'h149, 12'h14a, 12'h14a, 12'h14a, 12'h14b, 12'h14b, 12'h14b, 12'h14c, 12'h14c, 12'h14c, 12'h14d, 12'h14d, 12'h14d, 12'h14e, 12'h14e, 12'h14e, 12'h14f, 12'h14f, 12'h14f, 12'h150, 12'h150, 12'h150, 12'h151, 12'h151, 12'h151, 
12'h152, 12'h152, 12'h152, 12'h153, 12'h153, 12'h153, 12'h153, 12'h154, 12'h154, 12'h154, 12'h155, 12'h155, 12'h155, 12'h156, 12'h156, 12'h156, 12'h157, 12'h157, 12'h158, 12'h158, 12'h158, 12'h159, 12'h159, 12'h159, 12'h15a, 12'h15a, 12'h15a, 12'h15b, 12'h15b, 12'h15b, 12'h15c, 12'h15c, 12'h15c, 12'h15d, 12'h15d, 12'h15d, 12'h15e, 12'h15e, 12'h15e, 12'h15f, 12'h15f, 12'h15f, 12'h160, 12'h160, 12'h160, 12'h161, 12'h161, 12'h161, 12'h162, 12'h162, 12'h162, 12'h163, 12'h163, 12'h163, 12'h164, 12'h164, 12'h165, 12'h165, 12'h165, 12'h166, 12'h166, 12'h166, 12'h167, 12'h167, 12'h167, 12'h168, 12'h168, 12'h168, 12'h169, 12'h169, 12'h169, 12'h16a, 12'h16a, 12'h16a, 12'h16b, 12'h16b, 12'h16c, 12'h16c, 12'h16c, 12'h16d, 12'h16d, 12'h16d, 12'h16e, 12'h16e, 12'h16e, 12'h16f, 12'h16f, 12'h16f, 12'h170, 12'h170, 12'h171, 12'h171, 12'h171, 12'h172, 12'h172, 12'h172, 12'h173, 12'h173, 12'h173, 12'h174, 
12'h174, 12'h175, 12'h175, 12'h175, 12'h176, 12'h176, 12'h176, 12'h177, 12'h177, 12'h177, 12'h178, 12'h178, 12'h179, 12'h179, 12'h179, 12'h17a, 12'h17a, 12'h17a, 12'h17b, 12'h17b, 12'h17c, 12'h17c, 12'h17c, 12'h17d, 12'h17d, 12'h17d, 12'h17e, 12'h17e, 12'h17f, 12'h17f, 12'h17f, 12'h180, 12'h180, 12'h180, 12'h181, 12'h181, 12'h182, 12'h182, 12'h182, 12'h183, 12'h183, 12'h183, 12'h184, 12'h184, 12'h185, 12'h185, 12'h185, 12'h186, 12'h186, 12'h186, 12'h187, 12'h187, 12'h188, 12'h188, 12'h188, 12'h189, 12'h189, 12'h18a, 12'h18a, 12'h18a, 12'h18b, 12'h18b, 12'h18b, 12'h18c, 12'h18c, 12'h18d, 12'h18d, 12'h18d, 12'h18e, 12'h18e, 12'h18f, 12'h18f, 12'h18f, 12'h190, 12'h190, 12'h191, 12'h191, 12'h191, 12'h192, 12'h192, 12'h192, 12'h193, 12'h193, 12'h194, 12'h194, 12'h194, 12'h195, 12'h195, 12'h196, 12'h196, 12'h196, 12'h197, 12'h197, 12'h198, 12'h198, 12'h198, 12'h199, 12'h199, 12'h19a, 12'h19a, 
12'h19a, 12'h19b, 12'h19b, 12'h19c, 12'h19c, 12'h19c, 12'h19d, 12'h19d, 12'h19e, 12'h19e, 12'h19e, 12'h19f, 12'h19f, 12'h1a0, 12'h1a0, 12'h1a0, 12'h1a1, 12'h1a1, 12'h1a2, 12'h1a2, 12'h1a3, 12'h1a3, 12'h1a3, 12'h1a4, 12'h1a4, 12'h1a5, 12'h1a5, 12'h1a5, 12'h1a6, 12'h1a6, 12'h1a7, 12'h1a7, 12'h1a7, 12'h1a8, 12'h1a8, 12'h1a9, 12'h1a9, 12'h1aa, 12'h1aa, 12'h1aa, 12'h1ab, 12'h1ab, 12'h1ac, 12'h1ac, 12'h1ac, 12'h1ad, 12'h1ad, 12'h1ae, 12'h1ae, 12'h1af, 12'h1af, 12'h1af, 12'h1b0, 12'h1b0, 12'h1b1, 12'h1b1, 12'h1b2, 12'h1b2, 12'h1b2, 12'h1b3, 12'h1b3, 12'h1b4, 12'h1b4, 12'h1b4, 12'h1b5, 12'h1b5, 12'h1b6, 12'h1b6, 12'h1b7, 12'h1b7, 12'h1b7, 12'h1b8, 12'h1b8, 12'h1b9, 12'h1b9, 12'h1ba, 12'h1ba, 12'h1bb, 12'h1bb, 12'h1bb, 12'h1bc, 12'h1bc, 12'h1bd, 12'h1bd, 12'h1be, 12'h1be, 12'h1be, 12'h1bf, 12'h1bf, 12'h1c0, 12'h1c0, 12'h1c1, 12'h1c1, 12'h1c1, 12'h1c2, 12'h1c2, 12'h1c3, 12'h1c3, 12'h1c4, 12'h1c4, 
12'h1c5, 12'h1c5, 12'h1c5, 12'h1c6, 12'h1c6, 12'h1c7, 12'h1c7, 12'h1c8, 12'h1c8, 12'h1c9, 12'h1c9, 12'h1c9, 12'h1ca, 12'h1ca, 12'h1cb, 12'h1cb, 12'h1cc, 12'h1cc, 12'h1cd, 12'h1cd, 12'h1ce, 12'h1ce, 12'h1ce, 12'h1cf, 12'h1cf, 12'h1d0, 12'h1d0, 12'h1d1, 12'h1d1, 12'h1d2, 12'h1d2, 12'h1d2, 12'h1d3, 12'h1d3, 12'h1d4, 12'h1d4, 12'h1d5, 12'h1d5, 12'h1d6, 12'h1d6, 12'h1d7, 12'h1d7, 12'h1d8, 12'h1d8, 12'h1d8, 12'h1d9, 12'h1d9, 12'h1da, 12'h1da, 12'h1db, 12'h1db, 12'h1dc, 12'h1dc, 12'h1dd, 12'h1dd, 12'h1de, 12'h1de, 12'h1df, 12'h1df, 12'h1df, 12'h1e0, 12'h1e0, 12'h1e1, 12'h1e1, 12'h1e2, 12'h1e2, 12'h1e3, 12'h1e3, 12'h1e4, 12'h1e4, 12'h1e5, 12'h1e5, 12'h1e6, 12'h1e6, 12'h1e7, 12'h1e7, 12'h1e7, 12'h1e8, 12'h1e8, 12'h1e9, 12'h1e9, 12'h1ea, 12'h1ea, 12'h1eb, 12'h1eb, 12'h1ec, 12'h1ec, 12'h1ed, 12'h1ed, 12'h1ee, 12'h1ee, 12'h1ef, 12'h1ef, 12'h1f0, 12'h1f0, 12'h1f1, 12'h1f1, 12'h1f2, 12'h1f2, 12'h1f3, 
12'h1f3, 12'h1f4, 12'h1f4, 12'h1f5, 12'h1f5, 12'h1f5, 12'h1f6, 12'h1f6, 12'h1f7, 12'h1f7, 12'h1f8, 12'h1f8, 12'h1f9, 12'h1f9, 12'h1fa, 12'h1fa, 12'h1fb, 12'h1fb, 12'h1fc, 12'h1fc, 12'h1fd, 12'h1fd, 12'h1fe, 12'h1fe, 12'h1ff, 12'h1ff, 12'h200, 12'h200, 12'h201, 12'h201, 12'h202, 12'h202, 12'h203, 12'h203, 12'h204, 12'h204, 12'h205, 12'h205, 12'h206, 12'h206, 12'h207, 12'h207, 12'h208, 12'h208, 12'h209, 12'h209, 12'h20a, 12'h20b, 12'h20b, 12'h20c, 12'h20c, 12'h20d, 12'h20d, 12'h20e, 12'h20e, 12'h20f, 12'h20f, 12'h210, 12'h210, 12'h211, 12'h211, 12'h212, 12'h212, 12'h213, 12'h213, 12'h214, 12'h214, 12'h215, 12'h215, 12'h216, 12'h216, 12'h217, 12'h217, 12'h218, 12'h218, 12'h219, 12'h21a, 12'h21a, 12'h21b, 12'h21b, 12'h21c, 12'h21c, 12'h21d, 12'h21d, 12'h21e, 12'h21e, 12'h21f, 12'h21f, 12'h220, 12'h220, 12'h221, 12'h221, 12'h222, 12'h223, 12'h223, 12'h224, 12'h224, 12'h225, 12'h225, 12'h226, 
12'h226, 12'h227, 12'h227, 12'h228, 12'h228, 12'h229, 12'h22a, 12'h22a, 12'h22b, 12'h22b, 12'h22c, 12'h22c, 12'h22d, 12'h22d, 12'h22e, 12'h22e, 12'h22f, 12'h230, 12'h230, 12'h231, 12'h231, 12'h232, 12'h232, 12'h233, 12'h233, 12'h234, 12'h234, 12'h235, 12'h236, 12'h236, 12'h237, 12'h237, 12'h238, 12'h238, 12'h239, 12'h239, 12'h23a, 12'h23b, 12'h23b, 12'h23c, 12'h23c, 12'h23d, 12'h23d, 12'h23e, 12'h23e, 12'h23f, 12'h240, 12'h240, 12'h241, 12'h241, 12'h242, 12'h242, 12'h243, 12'h244, 12'h244, 12'h245, 12'h245, 12'h246, 12'h246, 12'h247, 12'h248, 12'h248, 12'h249, 12'h249, 12'h24a, 12'h24a, 12'h24b, 12'h24c, 12'h24c, 12'h24d, 12'h24d, 12'h24e, 12'h24e, 12'h24f, 12'h250, 12'h250, 12'h251, 12'h251, 12'h252, 12'h252, 12'h253, 12'h254, 12'h254, 12'h255, 12'h255, 12'h256, 12'h257, 12'h257, 12'h258, 12'h258, 12'h259, 12'h259, 12'h25a, 12'h25b, 12'h25b, 12'h25c, 12'h25c, 12'h25d, 12'h25e, 12'h25e, 
12'h25f, 12'h25f, 12'h260, 12'h261, 12'h261, 12'h262, 12'h262, 12'h263, 12'h264, 12'h264, 12'h265, 12'h265, 12'h266, 12'h267, 12'h267, 12'h268, 12'h268, 12'h269, 12'h26a, 12'h26a, 12'h26b, 12'h26b, 12'h26c, 12'h26d, 12'h26d, 12'h26e, 12'h26e, 12'h26f, 12'h270, 12'h270, 12'h271, 12'h271, 12'h272, 12'h273, 12'h273, 12'h274, 12'h275, 12'h275, 12'h276, 12'h276, 12'h277, 12'h278, 12'h278, 12'h279, 12'h279, 12'h27a, 12'h27b, 12'h27b, 12'h27c, 12'h27d, 12'h27d, 12'h27e, 12'h27e, 12'h27f, 12'h280, 12'h280, 12'h281, 12'h282, 12'h282, 12'h283, 12'h283, 12'h284, 12'h285, 12'h285, 12'h286, 12'h287, 12'h287, 12'h288, 12'h288, 12'h289, 12'h28a, 12'h28a, 12'h28b, 12'h28c, 12'h28c, 12'h28d, 12'h28e, 12'h28e, 12'h28f, 12'h28f, 12'h290, 12'h291, 12'h291, 12'h292, 12'h293, 12'h293, 12'h294, 12'h295, 12'h295, 12'h296, 12'h297, 12'h297, 12'h298, 12'h299, 12'h299, 12'h29a, 12'h29a, 12'h29b, 12'h29c, 12'h29c, 
12'h29d, 12'h29e, 12'h29e, 12'h29f, 12'h2a0, 12'h2a0, 12'h2a1, 12'h2a2, 12'h2a2, 12'h2a3, 12'h2a4, 12'h2a4, 12'h2a5, 12'h2a6, 12'h2a6, 12'h2a7, 12'h2a8, 12'h2a8, 12'h2a9, 12'h2aa, 12'h2aa, 12'h2ab, 12'h2ac, 12'h2ac, 12'h2ad, 12'h2ae, 12'h2ae, 12'h2af, 12'h2b0, 12'h2b0, 12'h2b1, 12'h2b2, 12'h2b2, 12'h2b3, 12'h2b4, 12'h2b4, 12'h2b5, 12'h2b6, 12'h2b6, 12'h2b7, 12'h2b8, 12'h2b8, 12'h2b9, 12'h2ba, 12'h2ba, 12'h2bb, 12'h2bc, 12'h2bd, 12'h2bd, 12'h2be, 12'h2bf, 12'h2bf, 12'h2c0, 12'h2c1, 12'h2c1, 12'h2c2, 12'h2c3, 12'h2c3, 12'h2c4, 12'h2c5, 12'h2c5, 12'h2c6, 12'h2c7, 12'h2c8, 12'h2c8, 12'h2c9, 12'h2ca, 12'h2ca, 12'h2cb, 12'h2cc, 12'h2cc, 12'h2cd, 12'h2ce, 12'h2cf, 12'h2cf, 12'h2d0, 12'h2d1, 12'h2d1, 12'h2d2, 12'h2d3, 12'h2d4, 12'h2d4, 12'h2d5, 12'h2d6, 12'h2d6, 12'h2d7, 12'h2d8, 12'h2d8, 12'h2d9, 12'h2da, 12'h2db, 12'h2db, 12'h2dc, 12'h2dd, 12'h2dd, 12'h2de, 12'h2df, 12'h2e0, 12'h2e0, 12'h2e1, 
12'h2e2, 12'h2e3, 12'h2e3, 12'h2e4, 12'h2e5, 12'h2e5, 12'h2e6, 12'h2e7, 12'h2e8, 12'h2e8, 12'h2e9, 12'h2ea, 12'h2ea, 12'h2eb, 12'h2ec, 12'h2ed, 12'h2ed, 12'h2ee, 12'h2ef, 12'h2f0, 12'h2f0, 12'h2f1, 12'h2f2, 12'h2f3, 12'h2f3, 12'h2f4, 12'h2f5, 12'h2f6, 12'h2f6, 12'h2f7, 12'h2f8, 12'h2f8, 12'h2f9, 12'h2fa, 12'h2fb, 12'h2fb, 12'h2fc, 12'h2fd, 12'h2fe, 12'h2fe, 12'h2ff, 12'h300, 12'h301, 12'h301, 12'h302, 12'h303, 12'h304, 12'h304, 12'h305, 12'h306, 12'h307, 12'h307, 12'h308, 12'h309, 12'h30a, 12'h30b, 12'h30b, 12'h30c, 12'h30d, 12'h30e, 12'h30e, 12'h30f, 12'h310, 12'h311, 12'h311, 12'h312, 12'h313, 12'h314, 12'h314, 12'h315, 12'h316, 12'h317, 12'h318, 12'h318, 12'h319, 12'h31a, 12'h31b, 12'h31b, 12'h31c, 12'h31d, 12'h31e, 12'h31f, 12'h31f, 12'h320, 12'h321, 12'h322, 12'h322, 12'h323, 12'h324, 12'h325, 12'h326, 12'h326, 12'h327, 12'h328, 12'h329, 12'h32a, 12'h32a, 12'h32b, 12'h32c, 12'h32d, 
12'h32e, 12'h32e, 12'h32f, 12'h330, 12'h331, 12'h332, 12'h332, 12'h333, 12'h334, 12'h335, 12'h336, 12'h336, 12'h337, 12'h338, 12'h339, 12'h33a, 12'h33a, 12'h33b, 12'h33c, 12'h33d, 12'h33e, 12'h33e, 12'h33f, 12'h340, 12'h341, 12'h342, 12'h342, 12'h343, 12'h344, 12'h345, 12'h346, 12'h347, 12'h347, 12'h348, 12'h349, 12'h34a, 12'h34b, 12'h34b, 12'h34c, 12'h34d, 12'h34e, 12'h34f, 12'h350, 12'h350, 12'h351, 12'h352, 12'h353, 12'h354, 12'h355, 12'h355, 12'h356, 12'h357, 12'h358, 12'h359, 12'h35a, 12'h35a, 12'h35b, 12'h35c, 12'h35d, 12'h35e, 12'h35f, 12'h35f, 12'h360, 12'h361, 12'h362, 12'h363, 12'h364, 12'h365, 12'h365, 12'h366, 12'h367, 12'h368, 12'h369, 12'h36a, 12'h36b, 12'h36b, 12'h36c, 12'h36d, 12'h36e, 12'h36f, 12'h370, 12'h371, 12'h371, 12'h372, 12'h373, 12'h374, 12'h375, 12'h376, 12'h377, 12'h377, 12'h378, 12'h379, 12'h37a, 12'h37b, 12'h37c, 12'h37d, 12'h37e, 12'h37e, 12'h37f, 12'h380, 
12'h381, 12'h382, 12'h383, 12'h384, 12'h385, 12'h385, 12'h386, 12'h387, 12'h388, 12'h389, 12'h38a, 12'h38b, 12'h38c, 12'h38c, 12'h38d, 12'h38e, 12'h38f, 12'h390, 12'h391, 12'h392, 12'h393, 12'h394, 12'h395, 12'h395, 12'h396, 12'h397, 12'h398, 12'h399, 12'h39a, 12'h39b, 12'h39c, 12'h39d, 12'h39e, 12'h39e, 12'h39f, 12'h3a0, 12'h3a1, 12'h3a2, 12'h3a3, 12'h3a4, 12'h3a5, 12'h3a6, 12'h3a7, 12'h3a8, 12'h3a8, 12'h3a9, 12'h3aa, 12'h3ab, 12'h3ac, 12'h3ad, 12'h3ae, 12'h3af, 12'h3b0, 12'h3b1, 12'h3b2, 12'h3b3, 12'h3b3, 12'h3b4, 12'h3b5, 12'h3b6, 12'h3b7, 12'h3b8, 12'h3b9, 12'h3ba, 12'h3bb, 12'h3bc, 12'h3bd, 12'h3be, 12'h3bf, 12'h3c0, 12'h3c1, 12'h3c1, 12'h3c2, 12'h3c3, 12'h3c4, 12'h3c5, 12'h3c6, 12'h3c7, 12'h3c8, 12'h3c9, 12'h3ca, 12'h3cb, 12'h3cc, 12'h3cd, 12'h3ce, 12'h3cf, 12'h3d0, 12'h3d1, 12'h3d2, 12'h3d3, 12'h3d3, 12'h3d4, 12'h3d5, 12'h3d6, 12'h3d7, 12'h3d8, 12'h3d9, 12'h3da, 12'h3db, 12'h3dc, 
12'h3dd, 12'h3de, 12'h3df, 12'h3e0, 12'h3e1, 12'h3e2, 12'h3e3, 12'h3e4, 12'h3e5, 12'h3e6, 12'h3e7, 12'h3e8, 12'h3e9, 12'h3ea, 12'h3eb, 12'h3ec, 12'h3ed, 12'h3ee, 12'h3ef, 12'h3f0, 12'h3f1, 12'h3f2, 12'h3f3, 12'h3f4, 12'h3f5, 12'h3f6, 12'h3f7, 12'h3f8, 12'h3f9, 12'h3fa, 12'h3fb, 12'h3fc, 12'h3fd, 12'h3fe, 12'h3ff, 12'h400};

//this function divides val by 2^10
    function [DWIDTH_IN+BITS-1:0] QUANTIZE_I;
        input [DWIDTH_IN-1:0] mval;
        begin
            QUANTIZE_I = mval * QUANT_VAL;
        end
    endfunction
/*
    function [DWIDTH_IN-1:0] DEQUANTIZE_I;
        input [DWIDTH_IN+BITS-1:0] mval;
        begin
            DEQUANTIZE_I = $floor(mval / QUANT_VAL);
        end
    endfunction

    function [DWIDTH_IN+BITS-1:0] QUANTIZE_F;
        input real mval;
        begin
            QUANTIZE_F = $floor(mval * (1.0 * QUANT_VAL)); //$floor converts to whole number(integer)
        end
    endfunction

    function real DEQUANTIZE_F;
        input [DWIDTH_IN+BITS-1:0] mval;
        begin
            DEQUANTIZE_F = $floor(mval / (1.0 * QUANT_VAL)); //$floor converts to whole number(integer)
        end
    endfunction
*/
//BRAM used for storing the input floating point data

    bram #(
        .BRAM_BUFFER_SIZE(IMG_SIZE),
        .BRAM_DATA_WIDTH(DWIDTH_IN),
        .BRAM_ADDR_WIDTH(BRAM_ADDR_WIDTH) //needs to match bram_addr_width
    ) my_mem( 
        .clock(clock),
        .reset(reset), //maybe change this to signal that goes high when new frame?
        .rd_addr(bram_addr),
        .wr_addr(bram_addr),
        .wr_en(bram_wr_en),
        .din(bram_din),
        .dout(bram_dout)
    );

    always @(posedge clock) begin
        if (reset == 1'b1) begin
            fifo_out_din <= 'b0;
            fifo_out_wr_en <= 1'b0;
            alpha <= 'b0;
            denominator <= 'b0;
            bram_addr <= 'b0;
            bram_wr_en <= 'b1;
            state <= PROLOGUE;
            move_on <= 1'b0;
            move_on2 <= 1'b0;
            exp_val <= 'b0;
        end else begin
            fifo_out_din <= fifo_out_din_c;
            fifo_out_wr_en <= fifo_out_wr_en_c;
            bram_addr <= bram_addr_c;
            bram_wr_en <= bram_wr_en;
            move_on <= move_on_c;
            move_on2 <= move_on2_c;
            alpha <= alpha_c;
            state <= next_state;
            denominator <= denominator_c;
            exp_val <= exp_val_c;
        end
    end

        //CAN USE A STATE MACHINE
        //State 0:
        //Write all of pixel data to bram until
        //we get to the end of the first image, 
        //and Get alpha
        //State 1:
        //iterate thru using lookup table to fill in values for out_imm 
        //and the denominator of the softmax func
        //State 2:
        //iterate thru all values in bram one more time using the 
        //denominator, and 
        //return denominator values to fifo_out_din
        

    
    always @* begin
        next_state = state;
        bram_addr_c = bram_addr;
        //bram_wr_en_c = bram_wr_en;
        bram_wr_en = 1'b0;
        bram_din = 'b0;
        denominator_c = denominator;
        alpha_c = alpha;
        fifo_in_rd_en = 1'b0;
        fifo_out_wr_en_c = 1'b0;
        fifo_out_din_c = 'b0;
        mval = 'b0;
        move_on_c = move_on;
        move_on2_c = move_on2;
        exp_val_c = exp_val;

        

        //converted_data = QUANTIZE_I(fifo_in_dout); //HERE TO DO: may need to quantize in values into fixed point(not sure, dont think I need to)

      
        case (state)
        //Read from fifo and find the alpha value
            PROLOGUE: begin
                
                //fill in values of exp table, and find 
                if (fifo_in_empty == 1'b0) begin
                    fifo_in_rd_en = 1'b1;

                    bram_addr_c = bram_addr + 1;
                    bram_wr_en = 1'b1;
                    bram_din = fifo_in_dout;

                    if (fifo_in_dout > alpha) begin //converted_data
                            alpha_c = fifo_in_dout; //converted_data
                    end
                    if (bram_addr == IMG_SIZE - 1) begin
                        move_on_c = 1'b1;
                        bram_addr_c = 'b0;
                        //next_state = MIDDLOGUE;

                    end 
                    //spend 1 cycle reading the first bram val so it is ready when we move onto middlogue
                    //I think we need to spend an extra cycle in this state to let bram catch up?
                    if(move_on == 1'b1) begin
                        bram_wr_en = 1'b0;
                        bram_addr_c = 'b0;
                        next_state = MIDDLOGUE;
                    end
                end 
            end

//potentially break up into 2 states:
//1 sets address 
//next one does all the calculations for mval etc.
            MIDDLOGUE: begin
                //if (fifo_in_empty == 1'b0 && fifo_out_full == 1'b0) begin

                //Don't read from fifo while we do this
                //also dont write to bram here
                //fifo_in_rd_en = 1'b0;
                bram_addr_c = bram_addr;
                bram_wr_en = 1'b0;

                next_state = BRAM_WR_STAGE;

                if(move_on2 == 1'b1) begin
                    next_state = EPILOGUE;
                end
                //Compute in[i] - alpha, and lookup that value in the table

                mval = (bram_dout - alpha);// & 12'hfff;

//WHEN ALPHA_VAL = BRAM_OUT, THIS DOES NOT RETRIEVE THE RIGHT VALUE
//should I change the value in the table at index 0? maybe...
                if (mval == 'b0) begin
                    exp_val_c = exp_arr[4096]; //if mval is alpha, then exp(0) = 1, which is 1024 quantized
                end else if ($signed(mval) < 32'shfffff000) begin
                    exp_val_c = 'b0;
                end else begin
                    exp_val_c = exp_arr[mval & 12'hfff];  //store exp_val back into bram somehow 
                end
                denominator_c = denominator + exp_val; //BRAM_DOUT will start ad address 0 in BRAM and continue on up
            end


            //state to let exp_val store into location in memory
            BRAM_WR_STAGE: begin
                bram_addr_c = bram_addr + 1;
                bram_wr_en = 1'b1;
                bram_din = exp_val;

                if (bram_addr == IMG_SIZE - 1) begin
                    move_on2_c = 1'b1;
                    bram_addr_c = 'b0;
                    fifo_out_wr_en_c = 1'b1;
                end
                next_state = MIDDLOGUE;
            end

            EPILOGUE: begin

                //TO DO: REPLACE DIVIDER WITH JULIAN'S DIVIDER MODULE
                if (fifo_out_full == 1'b0) begin
                    
                    fifo_out_wr_en_c = 1'b1;
                    fifo_out_din_c = QUANTIZE_I(bram_dout) / denominator; //QUANTIZE_I the bram_dout value
                    bram_addr_c = bram_addr + 1;

                    if (bram_addr >= IMG_SIZE-1) begin
                        next_state = TEMP_END_STATE;
                        bram_addr_c = 'b0;
                    end 
                end
            end

            TEMP_END_STATE: begin
                next_state = TEMP_END_STATE;
                //do nothing
                //todo: just go back to prologue from epilogue for new frame
            end
        endcase
    end 

endmodule
